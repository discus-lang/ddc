(* Top level module imports everything so that we have a
   nice make target to build the proofs. *)
Require Import DDC.Base.
Require Import DDC.Language.Simple.