(* Top level module imports everything so that we have a
   nice make target to build the proofs. *)
Require Import DDC.Base.

(* Simply Typed Lambda Calculus (STLC) *)
Require Import DDC.Language.Simple.

(* STLC with Fixpoints, Boolean choice and Naturals. *)
Require Import DDC.Language.SimplePCF.

(* STLC with mutable references. *)
Require Import DDC.Language.SimpleRef.

(* STLC with algebraic data types. *)
Require Import DDC.Language.SimpleData.

(* STLC with work and space resource types *)
Require Import DDC.Language.SimpleResource.

(* System-F. Like STLC, but with type abstraction and application. *)
Require Import DDC.Language.SystemF.

(* System-F2. Like System-F2 but with type-type application. *)
Require Import DDC.Language.SystemF2.

(* System-F2 with algebraic data types *)
Require Import DDC.Language.SystemF2Data.

(* System-F2 with algebraic data types and a mutable store. *)
Require Import DDC.Language.SystemF2Store.

(* System-F2 with region and effect types *)
Require Import DDC.Language.SystemF2Effect.